struct {
    
}